module picture_sender( );



endmodule
