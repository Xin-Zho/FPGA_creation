module data_trans_ethernet_control( 
    
);



endmodule
